`ifndef __MAPTABLE_V__
`define __MAPTABLE_V__

`timescale 1ns/100ps

module maptable(
  // Inputs
  input logic clock,
  input logic reset,
  input enable,
  input logic commit,
  input logic [4:0] rd_commit,
  input logic [`ROB_TAG_LEN-1:0] rob_entry_commit,
  input INST inst, //inst from decoding stage
  input logic [`ROB_TAG_LEN-1:0] rob_entry_in, // rob entry from ROB
  input logic [4:0] rd, // dest_reg from decoding stage
  input logic valid_wb, // valid from wb from ROB
  input logic [4:0] rd_wb, // dest_reg from wb
  input logic [`ROB_TAG_LEN-1:0] rob_entry_wb, // rob entry from wb from ROB
  input branch_pending,
  input kill, resolve,

  // Outputs
  output MAPTABLE_PACKET maptable_packet_rs1,
  output MAPTABLE_PACKET maptable_packet_rs2
);
  
  // Maptable and ready_tag
  logic [`ROB_TAG_LEN-1:0] maptable[31:0];
  logic ready_tag_table[31:0];

  logic [`ROB_TAG_LEN-1:0] maptable_buffer[31:0];
  logic ready_tag_table_buffer[31:0];


  // mapped rs1
  always_comb begin

    if (valid_wb && rob_entry_wb == maptable[inst.r.rs1]) begin
      // forwarding
      maptable_packet_rs1.rob_tag_ready = `TRUE;
    end
    else begin
      maptable_packet_rs1.rob_tag_ready = ready_tag_table[inst.r.rs1];
    end

    maptable_packet_rs1.rob_tag_val = maptable[inst.r.rs1];
  end

  // mapped rs2
  always_comb begin
    if (valid_wb && rob_entry_wb == maptable[inst.r.rs2]) begin
      // forwarding
      maptable_packet_rs2.rob_tag_ready = `TRUE;
    end
    else begin
      maptable_packet_rs2.rob_tag_ready = ready_tag_table[inst.r.rs2];
    end

    maptable_packet_rs2.rob_tag_val = maptable[inst.r.rs2];
  end

  always_ff @(posedge clock) begin
    if (reset) begin
      integer i;
      for (i = 0; i < 32; i++) begin
        maptable[i] = 0;
        ready_tag_table[i] = 0;
        maptable_buffer[i] = 0;
        ready_tag_table_buffer[i] = 0;
      end
    end

    if (resolve) begin
      maptable_buffer <= maptable;
      ready_tag_table_buffer <= ready_tag_table;
    end
    else if (kill) begin
      maptable <= maptable_buffer;
      ready_tag_table <= ready_tag_table_buffer;
    end

    if ((valid_wb) && (rd_wb != `ZERO_REG) && (rob_entry_wb == maptable[rd_wb])) begin
      ready_tag_table[rd_wb] = 1;
      if (!branch_pending) ready_tag_table_buffer[rd_wb] = 1;
    end
    if ((commit) && (rd_commit != `ZERO_REG) && (rob_entry_commit == maptable[rd_commit])) begin
      maptable[rd_commit] = 0;
      ready_tag_table[rd_commit] = 0;
      if (!branch_pending) begin
        maptable_buffer[rd_commit] = 0;
        ready_tag_table_buffer[rd_commit] = 0;
      end
    end
    if (enable && rd != `ZERO_REG) begin
      maptable[rd] = rob_entry_in;
      ready_tag_table[rd] = 0;
      if (!branch_pending) begin
        maptable_buffer[rd] = rob_entry_in;
        ready_tag_table_buffer[rd] = 0;
      end
    end
  end

endmodule
`endif
